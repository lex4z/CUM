`timescale 1ns / 1ps

module tb_lab102(
    
    );
    logic clk = 0;
    logic [31:0] din1;
    logic [31:0] din2;
    logic [31:0] dout;
    
    always #(5) clk = ~clk;
    
    lab102 test102(
        .clk(clk),
        .din1(din1),
        .din2(din2),
        .dout(dout)
    );
    
    initial begin
        // 0 10001010 11101000000000000000000
        // 1 10001110 00110101000000000000000
        
        //следует добавить проверку с бесконечностями
        
        din1 = 32'h42325604;
        din2 = 32'hC15AE76C;
        #10;
        
        din1 = 32'b01000011110001011001110000000000;
        din2 = 32'b01000100011111111000000000000000;
        #10;
        
        
        din1 = 32'b01000101011101000000000000000000;
        din2 = 32'b11000111000110101000000000000000;
        #10;
        
        din1 = 32'b11000011110001011000000000000000;
        din2 = 32'b01000100011111111000000000000000;
        #10;
        
        din1 = 32'b11000011110001011000000000000000;
        din2 = 32'b11000111000110101000000000000000;
        #10;
        
        din1 = 32'b11000011110001011000000000000000;
        din2 = 32'b01000011110001011000000000000000;
        #10;
        
        
        din1 = 32'b0;
        din2 = 32'b01000100011111111000000000000000;
        #10;
        
        din1 = 32'b01000100011111111000000000000000;
        din2 = 32'b0;
        #10;
        
        din1 = 32'b0;
        din2 = 32'b0;
        #10;
        
        
        $stop;
    end
endmodule
